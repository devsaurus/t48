-------------------------------------------------------------------------------
--
-- The Program Status Word (PSW).
-- Implements the PSW with its special bits.
--
-- All rights reserved
--
-------------------------------------------------------------------------------

configuration t48_psw_rtl_c0 of t48_psw is

  for rtl
  end for;

end t48_psw_rtl_c0;
