-------------------------------------------------------------------------------
--
-- The Conditional Branch Logic unit.
-- Decisions whether to take a jump or not are made here.
--
-- $Id: cond_branch-c.vhd,v 1.1 2004-03-23 21:24:33 arniml Exp $
--
-- Copyright (c) 2004, Arnim Laeuger (arniml@opencores.org)
--
-- All rights reserved
--
-------------------------------------------------------------------------------

configuration cond_branch_rtl_c0 of cond_branch is

  for rtl
  end for;

end cond_branch_rtl_c0;
