-------------------------------------------------------------------------------
--
-- T8243 Core
--
-- $Id: t8243_core-c.vhd,v 1.1 2006-07-13 22:53:56 arniml Exp $
--
-------------------------------------------------------------------------------

configuration t8243_core_rtl_c0 of t8243_core is

  for rtl
  end for;

end t8243_core_rtl_c0;
