-------------------------------------------------------------------------------
--
-- The Wishbone master module.
--
-- $Id: wb_master-c.vhd,v 1.1 2005-05-05 19:49:03 arniml Exp $
--
-- Copyright (c) 2004, Arnim Laeuger (arniml@opencores.org)
--
-- All rights reserved
--
-------------------------------------------------------------------------------

configuration wb_master_rtl_c0 of wb_master is

  for rtl
  end for;

end wb_master_rtl_c0;
