-------------------------------------------------------------------------------
--
-- The Timer/Counter unit.
--
-- $Id: timer-c.vhd,v 1.1 2004-03-23 21:31:53 arniml Exp $
--
-- All rights reserved
--
-------------------------------------------------------------------------------

configuration timer_rtl_c0 of timer is

  for rtl
  end for;

end timer_rtl_c0;
