-------------------------------------------------------------------------------
--
-- The Conditional Branch Logic unit.
-- Decisions whether to take a jump or not are made here.
--
-- $Id: cond_branch-c.vhd,v 1.2 2005-06-11 10:08:43 arniml Exp $
--
-- Copyright (c) 2004, Arnim Laeuger (arniml@opencores.org)
--
-- All rights reserved
--
-------------------------------------------------------------------------------

configuration t48_cond_branch_rtl_c0 of t48_cond_branch is

  for rtl
  end for;

end t48_cond_branch_rtl_c0;
