-------------------------------------------------------------------------------
--
-- $Id: dmem_ctrl_pack-p.vhd,v 1.1 2004-03-23 21:24:33 arniml Exp $
--
-- Copyright (c) 2004, Arnim Laeuger (arniml@opencores.org)
--
-- All rights reserved
--
-------------------------------------------------------------------------------

package dmem_ctrl_pack is

  -----------------------------------------------------------------------------
  -- Address Type Identifier
  -----------------------------------------------------------------------------
  type dmem_addr_ident_t is (DM_PLAIN,
                             DM_REG,
                             DM_STACK,
                             DM_STACK_HIGH);

end dmem_ctrl_pack;


-------------------------------------------------------------------------------
-- File History:
--
-- $Log: not supported by cvs2svn $
--
-------------------------------------------------------------------------------
