-------------------------------------------------------------------------------
--
-- The Interrupt Controller.
-- It collects the interrupt sources and notifies the decoder.
--
-- $Id: int-c.vhd,v 1.1 2004-03-23 21:31:52 arniml Exp $
--
-- All rights reserved
--
-------------------------------------------------------------------------------

configuration int_rtl_c0 of int is

  for rtl
  end for;

end int_rtl_c0;
