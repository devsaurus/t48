-------------------------------------------------------------------------------
--
-- The Program Status Word (PSW).
-- Implements the PSW with its special bits.
--
-- $Id: psw-c.vhd,v 1.1 2004-03-23 21:31:53 arniml Exp $
--
-- All rights reserved
--
-------------------------------------------------------------------------------

configuration psw_rtl_c0 of psw is

  for rtl
  end for;

end psw_rtl_c0;
