-------------------------------------------------------------------------------
--
-- The Timer/Counter unit.
--
-- $Id: timer-c.vhd,v 1.2 2005-06-11 10:08:43 arniml Exp $
--
-- All rights reserved
--
-------------------------------------------------------------------------------

configuration t48_timer_rtl_c0 of t48_timer is

  for rtl
  end for;

end t48_timer_rtl_c0;
