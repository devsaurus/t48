-------------------------------------------------------------------------------
--
-- $Id: clock_ctrl-c.vhd,v 1.1 2004-03-23 21:31:52 arniml Exp $
--
-- The clock control unit.
--
-------------------------------------------------------------------------------

configuration clock_ctrl_rtl_c0 of clock_ctrl is

  for rtl
  end for;

end clock_ctrl_rtl_c0;
