-------------------------------------------------------------------------------
--
-- The Interface Timing Checker.
--
-- $Id: if_timing-c.vhd,v 1.1 2004-04-25 16:24:10 arniml Exp $
--
-- Copyright (c) 2004, Arnim Laeuger (arniml@opencores.org)
--
-- All rights reserved
--
-------------------------------------------------------------------------------

configuration if_timing_behav_c0 of if_timing is

  for behav
  end for;

end if_timing_behav_c0;


-------------------------------------------------------------------------------
-- File History:
--
-- $Log: not supported by cvs2svn $
-------------------------------------------------------------------------------
