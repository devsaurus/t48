-------------------------------------------------------------------------------
--
-- $Id: t8048-c.vhd,v 1.1 2004-03-23 21:31:53 arniml Exp $
--
-------------------------------------------------------------------------------

configuration t8048_struct_c0 of t8048 is

  for struct

    for rom_1k_b : syn_rom
      use configuration work.syn_rom_altera_c0;
    end for;

    for ram_64_b : syn_ram
      use configuration work.syn_ram_altera_c0;
    end for;

    for t48_core_b : t48_core
      use configuration work.t48_core_struct_c0;
    end for;

  end for;

end t8048_struct_c0;
