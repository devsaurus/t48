-------------------------------------------------------------------------------
--
-- $Id$
--
-- The clock control unit.
--
-------------------------------------------------------------------------------

configuration t48_clock_ctrl_rtl_c0 of t48_clock_ctrl is

  for rtl
  end for;

end t48_clock_ctrl_rtl_c0;
