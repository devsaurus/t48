-------------------------------------------------------------------------------
--
-- The Program Memory control unit.
-- All operations related to the Program Memory are managed here.
--
-- $Id$
--
-- All rights reserved
--
-------------------------------------------------------------------------------

configuration t48_pmem_ctrl_rtl_c0 of t48_pmem_ctrl is

  for rtl
  end for;

end t48_pmem_ctrl_rtl_c0;
