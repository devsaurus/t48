-------------------------------------------------------------------------------
--
-- The Port 1 unit.
-- Implements the Port 1 logic.
--
-- $Id: p1-c.vhd,v 1.1 2004-03-23 21:31:52 arniml Exp $
--
-- All rights reserved
--
-------------------------------------------------------------------------------

configuration p1_rtl_c0 of p1 is

  for rtl
  end for;

end p1_rtl_c0;
