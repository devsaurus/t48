-------------------------------------------------------------------------------
--
-- $Id: t48_tb_pack-p.vhd,v 1.1 2004-03-23 21:24:33 arniml Exp $
--
-- Copyright (c) 2004, Arnim Laeuger (arniml@opencores.org)
--
-- All rights reserved
--
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

package t48_tb_pack is

  -- Accumulator visibilty
  signal tb_accu_s : std_logic_vector(7 downto 0);

end t48_tb_pack;
