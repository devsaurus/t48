-------------------------------------------------------------------------------
--
-- The Timer/Counter unit.
--
-- All rights reserved
--
-------------------------------------------------------------------------------

configuration t48_timer_rtl_c0 of t48_timer is

  for rtl
  end for;

end t48_timer_rtl_c0;
