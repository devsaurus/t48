-------------------------------------------------------------------------------
--
-- The Data Memory control unit.
-- All accesses to the Data Memory are managed here.
--
-- Copyright (c) 2004, Arnim Laeuger (arniml@opencores.org)
--
-- All rights reserved
--
-------------------------------------------------------------------------------

configuration t48_dmem_ctrl_rtl_c0 of t48_dmem_ctrl is

  for rtl
  end for;

end t48_dmem_ctrl_rtl_c0;
