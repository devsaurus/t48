-------------------------------------------------------------------------------
--
-- The T48 Bus Connector.
-- Multiplexes all drivers of the T48 bus.
--
-- $Id: bus_mux-c.vhd,v 1.2 2005-06-11 10:08:43 arniml Exp $
--
-- Copyright (c) 2004, Arnim Laeuger (arniml@opencores.org)
--
-- All rights reserved
--
-------------------------------------------------------------------------------

configuration t48_bus_mux_rtl_c0 of t48_bus_mux is

  for rtl
  end for;

end t48_bus_mux_rtl_c0;
