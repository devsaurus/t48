-------------------------------------------------------------------------------
--
-- The Opcode Decoder Table.
-- Decodes the given opcode to instruction mnemonics.
-- Also derives the multicycle information.
--
-- $Id: opc_table-c.vhd,v 1.1 2004-03-23 21:31:52 arniml Exp $
--
-- All rights reserved
--
-------------------------------------------------------------------------------

configuration opc_table_rtl_c0 of opc_table is

  for rtl
  end for;

end opc_table_rtl_c0;
