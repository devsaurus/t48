-------------------------------------------------------------------------------
--
-- The Program Memory control unit.
-- All operations related to the Program Memory are managed here.
--
-- $Id: pmem_ctrl-c.vhd,v 1.1 2004-03-23 21:24:33 arniml Exp $
--
-- All rights reserved
--
-------------------------------------------------------------------------------

configuration pmem_ctrl_rtl_c0 of pmem_ctrl is

  for rtl
  end for;

end pmem_ctrl_rtl_c0;
