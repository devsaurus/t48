-------------------------------------------------------------------------------
--
-- The Program Memory control unit.
-- All operations related to the Program Memory are managed here.
--
-- $Id: pmem_ctrl-c.vhd,v 1.2 2005-06-11 10:08:43 arniml Exp $
--
-- All rights reserved
--
-------------------------------------------------------------------------------

configuration t48_pmem_ctrl_rtl_c0 of t48_pmem_ctrl is

  for rtl
  end for;

end t48_pmem_ctrl_rtl_c0;
