-------------------------------------------------------------------------------
--
-- The Port 2 unit.
-- Implements the Port 2 logic.
--
-- $Id: p2.vhd,v 1.1 2004-03-23 21:24:33 arniml Exp $
--
-- All rights reserved
--
-- Redistribution and use in source and synthezised forms, with or without
-- modification, are permitted provided that the following conditions are met:
--
-- Redistributions of source code must retain the above copyright notice,
-- this list of conditions and the following disclaimer.
--
-- Redistributions in synthesized form must reproduce the above copyright
-- notice, this list of conditions and the following disclaimer in the
-- documentation and/or other materials provided with the distribution.
--
-- Neither the name of the author nor the names of other contributors may
-- be used to endorse or promote products derived from this software without
-- specific prior written permission.
--
-- THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS"
-- AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR
-- PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE AUTHOR OR CONTRIBUTORS BE
-- LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR
-- CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF
-- SUBSTITUTE GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS
-- INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN
-- CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE
-- POSSIBILITY OF SUCH DAMAGE.
--
-- Please report bugs to the author, but before you do so, please
-- make sure that this is not a derivative work and that
-- you have the latest version of this file.
--
-- The latest version of this file can be found at:
--      http://www.opencores.org/cvsweb.shtml/t48/
--
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

use work.t48_pack.word_t;
use work.t48_pack.nibble_t;

entity p2 is

  port (
    -- Global Interface -------------------------------------------------------
    clk_i        : in  std_logic;
    res_i        : in  std_logic;
    en_clk_i     : in  boolean;
    -- T48 Bus Interface ------------------------------------------------------
    data_i       : in  word_t;
    data_o       : out word_t;
    write_p2_i   : in  boolean;
    write_exp_i  : in  boolean;
    read_p2_i    : in  boolean;
    read_reg_i   : in  boolean;
    -- Port 2 Interface -------------------------------------------------------
    output_pch_i : in  boolean;
    output_exp_i : in  boolean;
    pch_i        : in  nibble_t;
    p2_i         : in  word_t;
    p2_o         : out word_t;
    p2_limp_o    : out std_logic
  );

end p2;


library ieee;
use ieee.std_logic_arith.conv_integer;
use ieee.std_logic_arith.unsigned;

use work.t48_pack.clk_active_c;
use work.t48_pack.res_active_c;
use work.t48_pack.bus_idle_level_c;

architecture rtl of p2 is

  subtype exp_t  is std_logic_vector(1 downto 0);

  -- 8243 expander address mapping
  type     exp_array_t is array (3 downto 0) of nibble_t;
  constant exp_c : exp_array_t := ("0100", "0101", "0110", "0111");

  -- the port output register
  signal p2_q   : word_t;

  -- the low impedance marker
  signal limp_q : std_logic;

  -- the expander register
  signal exp_q  : exp_t;
  signal exp_s  : nibble_t;

begin

  -----------------------------------------------------------------------------
  -- Process p2_regs
  --
  -- Purpose:
  --   Implements the port output and expander registers.
  --
  p2_regs: process (res_i, clk_i)
  begin
    if res_i = res_active_c then
      p2_q     <= (others => '1');
      limp_q   <= '0';
      exp_q    <= (others => '0');

    elsif clk_i'event and clk_i = clk_active_c then
      if en_clk_i then

        if write_p2_i then
          p2_q   <= data_i;
          limp_q <= '1';
        else
          limp_q <= '0';
        end if;

        if write_exp_i then
          exp_q  <= data_i(exp_q'range);
        end if;

      end if;

    end if;

  end process p2_regs;
  --
  -----------------------------------------------------------------------------


  exp_s <= exp_c(conv_integer(unsigned(exp_q)));


  -----------------------------------------------------------------------------
  -- Output Mapping.
  -----------------------------------------------------------------------------
  p2_o      <=   "0000" & exp_s
               when output_exp_i else
                 "0000" & pch_i
               when output_pch_i else
                 p2_q;
  p2_limp_o <= limp_q;

  data_o    <=   (others => bus_idle_level_c)
               when not read_p2_i else
                 p2_q
               when read_reg_i else
                 p2_i;

end rtl;


-------------------------------------------------------------------------------
-- File History:
--
-- $Log: not supported by cvs2svn $
--
-------------------------------------------------------------------------------
