-------------------------------------------------------------------------------
--
-- The Interrupt Controller.
-- It collects the interrupt sources and notifies the decoder.
--
-- $Id$
--
-- All rights reserved
--
-------------------------------------------------------------------------------

configuration t48_int_rtl_c0 of t48_int is

  for rtl
  end for;

end t48_int_rtl_c0;
