-------------------------------------------------------------------------------
--
-- The Interrupt Controller.
-- It collects the interrupt sources and notifies the decoder.
--
-- $Id: int-c.vhd,v 1.2 2005-06-11 10:08:43 arniml Exp $
--
-- All rights reserved
--
-------------------------------------------------------------------------------

configuration t48_int_rtl_c0 of t48_int is

  for rtl
  end for;

end t48_int_rtl_c0;
