-------------------------------------------------------------------------------
--
-- The T48 Bus Connector.
-- Multiplexes all drivers of the T48 bus.
--
-- Copyright (c) 2004, Arnim Laeuger (arniml@opencores.org)
--
-- All rights reserved
--
-------------------------------------------------------------------------------

configuration t48_bus_mux_rtl_c0 of t48_bus_mux is

  for rtl
  end for;

end t48_bus_mux_rtl_c0;
