-------------------------------------------------------------------------------
--
-- T8243 Core
--
-- $Id$
--
-------------------------------------------------------------------------------

configuration t8243_core_rtl_c0 of t8243_core is

  for rtl
  end for;

end t8243_core_rtl_c0;
