-------------------------------------------------------------------------------
--
-- The Port 2 unit.
-- Implements the Port 2 logic.
--
-- All rights reserved
--
-------------------------------------------------------------------------------

configuration t48_p2_rtl_c0 of t48_p2 is

  for rtl
  end for;

end t48_p2_rtl_c0;
