-------------------------------------------------------------------------------
--
-- The Interface Timing Checker.
--
-- Copyright (c) 2004, Arnim Laeuger (arniml@opencores.org)
--
-- All rights reserved
--
-------------------------------------------------------------------------------

configuration if_timing_behav_c0 of if_timing is

  for behav
  end for;

end if_timing_behav_c0;
