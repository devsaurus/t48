-------------------------------------------------------------------------------
--
-- The T48 SAR ADC.
--
-- Copyright (c) 2023, Arnim Laeuger (arniml@opencores.org)
--
-- All rights reserved
--
-------------------------------------------------------------------------------

configuration t48_adc_rtl_c0 of t48_adc is

  for rtl
  end for;

end t48_adc_rtl_c0;
