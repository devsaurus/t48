-------------------------------------------------------------------------------
--
-- The BUS unit.
-- Implements the BUS port logic.
--
-- Copyright (c) 2004, Arnim Laeuger (arniml@opencores.org)
--
-- All rights reserved
--
-------------------------------------------------------------------------------

configuration t48_db_bus_rtl_c0 of t48_db_bus is

  for rtl
  end for;

end t48_db_bus_rtl_c0;
