-------------------------------------------------------------------------------
--
-- The Port 1 unit.
-- Implements the Port 1 logic.
--
-- $Id$
--
-- All rights reserved
--
-------------------------------------------------------------------------------

configuration t48_p1_rtl_c0 of t48_p1 is

  for rtl
  end for;

end t48_p1_rtl_c0;
