-------------------------------------------------------------------------------
--
-- The Data Memory control unit.
-- All accesses to the Data Memory are managed here.
--
-- $Id: dmem_ctrl-c.vhd,v 1.1 2004-03-23 21:31:52 arniml Exp $
--
-- Copyright (c) 2004, Arnim Laeuger (arniml@opencores.org)
--
-- All rights reserved
--
-------------------------------------------------------------------------------

configuration dmem_ctrl_rtl_c0 of dmem_ctrl is

  for rtl
  end for;

end dmem_ctrl_rtl_c0;
