
configuration upi_stim_behav_c0 of upi_stim is

  for behav
  end for;

end upi_stim_behav_c0;
