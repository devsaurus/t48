-------------------------------------------------------------------------------
--
-- The Port 2 unit.
-- Implements the Port 2 logic.
--
-- $Id: p2-c.vhd,v 1.1 2004-03-23 21:31:53 arniml Exp $
--
-- All rights reserved
--
-------------------------------------------------------------------------------

configuration p2_rtl_c0 of p2 is

  for rtl
  end for;

end p2_rtl_c0;
